`timescale 1ns/1ps;
module accumulation_32_tb;
reg clk;
reg rstn;
reg en;
wire done;
reg [255:0] feature;
reg [255:0] weight;
wire [19:0] result;
reg signed [19:0] partial_sum [0:7];
reg signed [20:0] tmp_adder4 [0:3];
reg signed [21:0] tmp_adder2 [0:1];
reg signed [22:0] tmp_adder1;
reg signed [7:0] bias;
reg [3:0] iter;
reg [7:0] out;
integer i;

parameter CLK_CYCLE = 5;

accumulation_32 dut (
    .clk(clk),
    .rstn(rstn),
    .en(en),
    .done(done),
    .feature(feature),
    .weight(weight),
    .result(result)
);

always #CLK_CYCLE clk = ~clk;

initial begin
    clk = 1'b0;
    rstn = 1'b0;
    en = 1'b0;
    iter = 4'b0;
    bias = {8{1'b0}};
    tmp_adder4[0] = {21{1'b0}};
    tmp_adder4[1] = {21{1'b0}};
    tmp_adder4[2] = {21{1'b0}};
    tmp_adder4[3] = {21{1'b0}};
    tmp_adder2[0] = {22{1'b0}};
    tmp_adder2[1] = {22{1'b0}};
    tmp_adder1 = {23{1'b0}};

    for (i = 0; i < 8; i = i + 1) begin
        partial_sum[i] = {20{1'b0}};
    end

    repeat(5)
        @(posedge clk)

    rstn = 1'b1;

    repeat(5)
        @(posedge clk)

    feature[31:0]    = 32'b00010000000011110001110100000000;
    feature[63:32]   = 32'b00001101000001100000000000000000;
    feature[95:64]   = 32'b00000000000011110000100100011101;
    feature[127:96]  = 32'b00000000000000000000000100001101;
    feature[159:128] = 32'b00000001000001000000011000000000;
    feature[191:160] = 32'b00010001000011010001000100000011;
    feature[223:192] = 32'b00010111000111100000000000001101;
    feature[255:224] = 32'b00001111000110110010011000001110;

    weight[31:0]     = 32'b00000000000000001111110100000000;
    weight[63:32]    = 32'b11111101111111100000000000000000;
    weight[95:64]    = 32'b00000001000000000000000100001001;
    weight[127:96]   = 32'b00000000000000000000000111111110;
    weight[159:128]  = 32'b00000001000000001111110000000000;
    weight[191:160]  = 32'b00000000111111111111111100000010;
    weight[223:192]  = 32'b11111000111111010000001111111111;
    weight[255:224]  = 32'b11111010000000010000011100000010;

    repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = iter + 4'b1;
    en = 1'b0;

    repeat(5)
        @(posedge clk)
    
    // ft - I_63
    feature[31:0]    = 32'b00010001000010000000111000000000;
    feature[63:32]   = 32'b00010111000000010000100000001011;
    feature[95:64]   = 32'b00000000000100100001101000010000;
    feature[127:96]  = 32'b00000111000011000000000000011110;
    feature[159:128] = 32'b00001100000101000000011100010010;
    feature[191:160] = 32'b00001100000100100000000000000100;
    feature[223:192] = 32'b00010000000000000000000000000111;
    feature[255:224] = 32'b00000000000000100000101100000001;


    // wt - W_63
    weight[31:0]     = 32'b00000000000000000000000111111111;
    weight[63:32]    = 32'b00000000111111110000010100000010;
    weight[95:64]    = 32'b00000000111110101111100100000100;
    weight[127:96]   = 32'b00000011111111100000000011111110;
    weight[159:128]  = 32'b11111110000000000000000000000000;
    weight[191:160]  = 32'b11111110111111000000000000000001;
    weight[223:192]  = 32'b00000010000000000000000000000001;
    weight[255:224]  = 32'b00000000000000000000000000000001;

    repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = iter + 4'b1;
    en = 1'b0;

    repeat(5)
        @(posedge clk)

    // ft - I _95
    feature[31:0]    = 32'b00001111000011000000000000010000;
    feature[63:32]   = 32'b00001010000000000000111000100000;
    feature[95:64]   = 32'b00011000000011110001100000010100;
    feature[127:96]  = 32'b00010000000000000000110000000111;
    feature[159:128] = 32'b00000111000000000001010000000000;
    feature[191:160] = 32'b00000000000000000000000000000101;
    feature[223:192] = 32'b00011011000000000000111100000000;
    feature[255:224] = 32'b00000000000000000001000000000111;

    // wt - W_95
    weight[31:0]     = 32'b00010001000010000000111000000000;
    weight[63:32]    = 32'b00010111000000010000100000001011;
    weight[95:64]    = 32'b00000000000100100001101000010000;
    weight[127:96]   = 32'b00000111000011000000000000011110;
    weight[159:128]  = 32'b00001100000101000000011100010010;
    weight[191:160]  = 32'b00001100000100100000000000000100;
    weight[223:192]  = 32'b00010000000000000000000000000111;
    weight[255:224]  = 32'b00000000000000100000101100000001;

    repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = iter + 4'b1;
    en = 1'b0;

    repeat(5)
        @(posedge clk)

    // ft - I _127
    feature[31:0]    = 32'b00001110000010010000000000010111;
    feature[63:32]   = 32'b00000000000101110001101000011110;
    feature[95:64]   = 32'b00000000000100010001001000011100;
    feature[127:96]  = 32'b00000010000111000000011100000011;
    feature[159:128] = 32'b00000000000001000000000000010000;
    feature[191:160] = 32'b00001101000101010001100000000000;
    feature[223:192] = 32'b00001010000010100001000000000000;
    feature[255:224] = 32'b00001010000000000000101000010011;

    // wt - W_127
    weight[31:0]     = 32'b11111110000001000000000000010000;
    weight[63:32]    = 32'b00000000000000000000001111111100;
    weight[95:64]    = 32'b00000000000001010000100011111010;
    weight[127:96]   = 32'b00000010111110110000000011111111;
    weight[159:128]  = 32'b00000000111111110000000000000011;
    weight[191:160]  = 32'b00000000000000100000111000000000;
    weight[223:192]  = 32'b11111111111111011111110100000000;
    weight[255:224]  = 32'b11111110000000000000100011111101;

    repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = iter + 4'b1;
    en = 1'b0;

    repeat(5)
        @(posedge clk)

    // ft - I _159
    feature[31:0]    = 32'b00001110000101100000100100000000;
    feature[63:32]   = 32'b00000101000001100000100100100000;
    feature[95:64]   = 32'b00000000000000000000101000000010;
    feature[127:96]  = 32'b00001110000000100000000000000000;
    feature[159:128] = 32'b00010001000010000000001000001001;
    feature[191:160] = 32'b00000000000011100000111000001111;
    feature[223:192] = 32'b00000110000000110001000100000000;
    feature[255:224] = 32'b00000000000000110001010100001111;

    // wt - W_159
    weight[31:0]     = 32'b00000100000100001111110100000000;
    weight[63:32]    = 32'b00000000111110100000010100000000;
    weight[95:64]    = 32'b00000000000000001111111111111111;
    weight[127:96]   = 32'b00000000000000110000000000000000;
    weight[159:128]  = 32'b00000000111111100000000000000000;
    weight[191:160]  = 32'b00000000000000111111110111111111;
    weight[223:192]  = 32'b00000011000000000000001000000000;
    weight[255:224]  = 32'b00000000000000000000101111111101;
    
     repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = iter + 4'b1;
    en = 1'b0;

    repeat(5)
        @(posedge clk)

    // ft - I _191
    feature[31:0]    = 32'b00001110000000000001001100000000;
    feature[63:32]   = 32'b00000000000100010001001000001110;
    feature[95:64]   = 32'b00000101000011100001010000000011;
    feature[127:96]  = 32'b00000000000000000000100100000000;
    feature[159:128] = 32'b00000000000011010000100100011010;
    feature[191:160] = 32'b00001101000101110000000000000001;
    feature[223:192] = 32'b00000000000010010001010000000000;
    feature[255:224] = 32'b00000000000110010000011000001001;

    // wt - W_191
    weight[31:0]     = 32'b00000011000000001111101100000000;
    weight[63:32]    = 32'b00000000000000000000001000000100;
    weight[95:64]    = 32'b00000010111110011111100000000011;
    weight[127:96]   = 32'b00000000000000000000010000000000;
    weight[159:128]  = 32'b00000000000000001111111100001001;
    weight[191:160]  = 32'b00000000111110110000000000000001;
    weight[223:192]  = 32'b00000000000001100000010000000000;
    weight[255:224]  = 32'b00000000111111000000000011111011;

    repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = iter + 4'b1;
    en = 1'b0;

    repeat(5)
        @(posedge clk)

    // ft - I _223
    feature[31:0]    = 32'b00000110001000110000000000000000;
    feature[63:32]   = 32'b00000000000000000000111100000000;
    feature[95:64]   = 32'b00011100000010100000000000000100;
    feature[127:96]  = 32'b00001010000000000000000000000011;
    feature[159:128] = 32'b00000101001011000000000000001000;
    feature[191:160] = 32'b00001101000100000000101100000111;
    feature[223:192] = 32'b00000000000011010000000000000010;
    feature[255:224] = 32'b00001111000010110000111000001100;

    // wt - W_223
    weight[31:0]     = 32'b00000001111111010000000000000000;
    weight[63:32]    = 32'b00000000000000000000010000000000;
    weight[95:64]    = 32'b11111110000000000000000000000001;
    weight[127:96]   = 32'b00000110000000000000000000000001;
    weight[159:128]  = 32'b00000000000001000000000000000011;
    weight[191:160]  = 32'b11111010111111100000000000000110;
    weight[223:192]  = 32'b00000000000000000000000000000000;
    weight[255:224]  = 32'b00000000000000100000000100000001;

    repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = iter + 4'b1;
    en = 1'b0;

    repeat(5)
        @(posedge clk)

    // ft - I _255
    feature[31:0]    = 32'b00000000000010110001100100001001;
    feature[63:32]   = 32'b00000000000100100001000100000000;
    feature[95:64]   = 32'b00010011000111110000000000000111;
    feature[127:96]  = 32'b00000000000001100001100100000010;
    feature[159:128] = 32'b00000000000000000000000000000000;
    feature[191:160] = 32'b00000000000100100000000100000000;
    feature[223:192] = 32'b00010011000000000000110100010100;
    feature[255:224] = 32'b00001001000100110000101000011011;

    // wt - W_255
    weight[31:0]     = 32'b00000000000000000000001000000100;
    weight[63:32]    = 32'b00000000000101010000001100000000;
    weight[95:64]    = 32'b00000001000001000000000000000000;
    weight[127:96]   = 32'b00000001111111110001000000000000;
    weight[159:128]  = 32'b00000000000000000000000000000000;
    weight[191:160]  = 32'b00000000000010000000000000000000;
    weight[223:192]  = 32'b11111111000000001111110100000000;
    weight[255:224]  = 32'b00000001000000000000100000001011;

    repeat(5)
        @(posedge clk)
    en = 1'b1;

    wait(done)
    $display("The partial sum is: %b", result);
    partial_sum[iter] = result;
    iter = 4'b0;
    en = 1'b0;

    repeat(5)
        @(posedge clk)

    tmp_adder4[0] = partial_sum[0] + partial_sum[1];
    tmp_adder4[1] = partial_sum[2] + partial_sum[3];
    tmp_adder4[2] = partial_sum[4] + partial_sum[5];
    tmp_adder4[3] = partial_sum[6] + partial_sum[7];

    repeat(5)
        @(posedge clk)

    tmp_adder2[0] = tmp_adder4[0] + tmp_adder4[1];
    tmp_adder2[1] = tmp_adder4[2] + tmp_adder4[3];

    repeat(5)
        @(posedge clk)

    tmp_adder1 = tmp_adder2[0] + tmp_adder2[1] + bias;

    repeat(5)
        @(posedge clk)

    $display("tmp_adder1_value: %b", tmp_adder1);
    // qunatization
    if (tmp_adder1[21:13] == {9{1'b0}} || tmp_adder1[21:13] == {9{1'b1}}) begin
        out[7] = tmp_adder1[22];
        out[6:0] = tmp_adder1[12:6];
    end
    else if (tmp_adder1[22] == 1'b1) begin
    // negative OF
        out = 8'b1000_0000;
    end
    else begin
    // positive OF
        out = 8'b0111_1111;
    end

    repeat(5)
        @(posedge clk)

    // relu
    if (out[7] == 1'b1) out = 8'b0000_0000;

    $display("The output value is: %b", out);

    $finish;
end

endmodule